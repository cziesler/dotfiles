module hello_world();

initial begin
  $display ("Hello, world!");
end

endmodule
